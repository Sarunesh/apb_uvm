interface apb_intf(input logic pclk, input logic preset_n);
endinterface
