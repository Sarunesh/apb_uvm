`include "uvm_pkg.sv"
import uvm_pkg::*;
`include "apb.v"
`include "mem.v"
`include "apb_common.sv"
`include "apb_intf.sv"
`include "apb_tx.sv"
`include "apb_seq_lib.sv"
`include "apb_sqr.sv"
`include "apb_drv.sv"
`include "apb_mon.sv"
`include "apb_sub.sv"
`include "apb_agent.sv"
`include "apb_sbd.sv"
`include "apb_env.sv"
`include "test_lib.sv"
`include "top.sv"
