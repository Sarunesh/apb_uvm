class apb_seq_lib extends uvm_sequence#(apb_tx);
	// Factory registration
	`uvm_object_utils(apb_seq_lib)

	// Constructor
	`NEW_OBJECT
endclass
