class apb_tx extends uvm_sequence_item;
	// Properties

	// Factory registration
	`uvm_object_utils_begin(apb_tx)
	`uvm_object_utils_end

	// Constructor
	`NEW_OBJECT
endclass
